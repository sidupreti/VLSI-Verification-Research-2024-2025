module Benchmarks/2n+1/4( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31_0 , n31_1 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39_0 , n39_1 , n40 , n41_0 , n41_1 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53_0 , n53_1 , n54 , n55_0 , n55_1 , n56_0 , n56_1 , n57 , n58 , n59 , n60_0 , n60_1 , n61 , n62_0 , n62_1 , n63 , n64_0 , n64_1 , n65 , n67_0 , n67_1 , n68 , n70_0 , n70_1 ;
  AND               g00( .A (x2), .B (x5), .Y (n21) );
  INV               g01( .A (n21), .Y (n22) );
  AND               g02( .A (x3), .B (x4), .Y (n23) );
  INV               g03( .A (n23), .Y (n24) );
  AND               g04( .A (x0), .B (x7), .Y (n25) );
  INV               g05( .A (n25), .Y (n26) );
  AND               g06( .A (n24), .B (n26), .Y (n27) );
  AND               g07( .A (n22), .B (n27), .Y (n28) );
  INV               g08( .A (n28), .Y (n29) );
  AND               g09( .A (x1), .B (x6), .Y (n30) );
  AND               g10( .A (x3), .B (x7), .Y (n18) );
  INV               g11( .A (n18), .Y (n19) );
  AND               g12( .A (x0), .B (x4), .Y (n10) );
  INV               g13( .A (n10), .Y (n11) );
  AND               g14( .A (x3), .B (x6), .Y (n12) );
  INV               g15( .A (n12), .Y (n13) );
  AND               g16( .A (x2), .B (x7), .Y (n14) );
  INV               g17( .A (n14), .Y (n15) );
  AND               g18( .A (n13), .B (n15), .Y (n16) );
  AND               g19( .A (n11), .B (n16), .Y (n17) );
  AND               g20( .A (n19), .B (n17), .Y (n20) );
  FA                g21( .A (n29), .B (n30), .CI (n20), .CON (n31_0), .SN (n31_1) );
  AND               g22( .A (x2), .B (x4), .Y (n35) );
  INV               g23( .A (n35), .Y (n36) );
  AND               g24( .A (n36), .B (n16), .Y (n37) );
  INV               g25( .A (n37), .Y (n38) );
  AND               g26( .A (x1), .B (x5), .Y (n34) );
  AND               g27( .A (x0), .B (x6), .Y (n33) );
  FA                g28( .A (n38), .B (n34), .CI (n33), .CON (n39_0), .SN (n39_1) );
  HA                g29( .A (n31_1), .B (n39_0), .CON (n41_0), .SN (n41_1) );
  INV               g30( .A (n41_1), .Y (n42) );
  AND               g31( .A (x0), .B (x5), .Y (n43) );
  AND               g32( .A (x1), .B (x4), .Y (n44) );
  AND               g33( .A (x2), .B (x6), .Y (n45) );
  INV               g34( .A (n45), .Y (n46) );
  AND               g35( .A (x3), .B (x5), .Y (n47) );
  INV               g36( .A (n47), .Y (n48) );
  AND               g37( .A (x1), .B (x7), .Y (n49) );
  INV               g38( .A (n49), .Y (n50) );
  AND               g39( .A (n48), .B (n50), .Y (n51) );
  AND               g40( .A (n46), .B (n51), .Y (n52) );
  FA                g41( .A (n43), .B (n44), .CI (n52), .CON (n53_0), .SN (n53_1) );
  INV               g42( .A (n53_0), .Y (n54) );
  INV               g43( .A (n39_1), .Y (n40) );
  HA                g44( .A (n54), .B (n40), .CON (n55_0), .SN (n55_1) );
  HA                g45( .A (n42), .B (n55_0), .CON (n56_0), .SN (n56_1) );
  INV               g46( .A (n56_1), .Y (n57) );
  INV               g47( .A (n31_0), .Y (n32) );
  AND               g48( .A (n32), .B (n53_1), .Y (n59) );
  XOR               g49( .A (n32), .B (n53_1), .Y (n58) );
  FA                g50( .A (n41_0), .B (n56_0), .CI (n58), .CON (n60_0), .SN (n60_1) );
  INV               g51( .A (n60_0), .Y (n61) );
  FA                g52( .A (n59), .B (n55_1), .CI (n61), .CON (n62_0), .SN (n62_1) );
  INV               g53( .A (n62_0), .Y (n63) );
  HA                g54( .A (n57), .B (n63), .CON (n64_0), .SN (n64_1) );
  INV               g55( .A (n64_1), .Y (y0) );
  INV               g56( .A (n64_0), .Y (n65) );
  HA                g57( .A (n60_1), .B (n65), .CON (n67_0), .SN (n67_1) );
  INV               g58( .A (n67_1), .Y (y1) );
  INV               g59( .A (n67_0), .Y (n68) );
  HA                g60( .A (n62_1), .B (n68), .CON (n70_0), .SN (n70_1) );
  INV               g61( .A (n70_1), .Y (y2) );
  INV               g62( .A (n70_0), .Y (y3) );
endmodule
